/**
    File: CoreDatapath.v
    Author: BlackIsDevin (https://github.com/BlackIsDevin)
    Date: 6/30/2021
    Target Devices:
        Mimas A7 Revision V3 Development Board
        Arty A7-35T Development Board (future target)
    Description:
        This modules holds the central datapath of the CPU core, as well as
        exposes parts of data memory (and in the future, a writable instruction
        memory module) to other modules.
*/


module CoreDatapath(
    input clk
);
    // TODO: literally all of this
endmodule
