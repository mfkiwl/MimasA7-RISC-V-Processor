// this modules holds the central datapath of the CPU core, as well as exposes 
// parts of data memory (and in the future, a writable instruction memory
// module) to other modules
module CoreDatapath(

);
    // TODO: literally all of this
endmodule