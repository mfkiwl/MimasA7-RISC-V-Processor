/**
    This modules holds the central datapath of the CPU core, as well as
        exposes parts of data memory (and in the future, a writable instruction
        memory module) to other modules.
    @author BlackIsDevin (https://github.com/BlackIsDevin)
    
        
*/


module CoreDatapath(
    input clk
);
    // TODO: literally all of this
endmodule
